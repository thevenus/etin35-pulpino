/usr/local-eit/cad2/cmpstm/oldmems/mem2010/SPHDL100909-40446@1.0/CADENCE/LEF/SPHDL100909_soc.lef