-- Top module for apb_conv connecting controller and convolve unit 