-- Convolution controller design